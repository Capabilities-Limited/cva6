// Copyright 2018 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

// Xilinx Peripherals

`include "register_interface/assign.svh"
`include "register_interface/typedef.svh"

module ariane_peripherals #(
    parameter int AxiAddrWidth = -1,
    parameter int AxiDataWidth = -1,
    parameter int AxiIdWidth   = -1,
    parameter int AxiUserWidth = 1,
    parameter bit InclUART     = 1,
    parameter bit InclSPI      = 0,
    parameter bit InclXilinxEthernet  = 0,
    parameter bit InclLowriscEthernet = 0,
    parameter bit InclGPIO     = 0,
    parameter bit InclTimer    = 1
) (
    input  logic       clk_i           , // Clock
    input  logic       clk_200MHz_i    ,
    input  logic       rst_ni          , // Asynchronous reset active low
    AXI_BUS.Slave      plic            ,
    AXI_BUS.Slave      uart            ,
    AXI_BUS.Slave      spi             ,
    AXI_BUS.Slave      gpio            ,
    AXI_BUS.Slave      ethernet_mgmt   ,
    AXI_BUS.Slave      ethernet_data   ,
    AXI_BUS.Slave      timer           ,
    output logic [1:0] irq_o           ,
    // UART
    input  logic       rx_i            ,
    output logic       tx_o            ,
    // Ethernet
    input  logic       eth_clk_i       ,
    input  wire        eth_rxck        ,
    input  wire        eth_rxctl       ,
    input  wire [3:0]  eth_rxd         ,
    output wire        eth_txck        ,
    output wire        eth_txctl       ,
    output wire [3:0]  eth_txd         ,
    output wire        eth_rst_n       ,
    input  logic       phy_tx_clk_i    , // 125 MHz Clock
    // MDIO Interface
    inout  wire        eth_mdio        ,
    output logic       eth_mdc         ,
    // SPI
    output logic       spi_clk_o       ,
    output logic       spi_mosi        ,
    input  logic       spi_miso        ,
    output logic       spi_ss          ,
    // SD Card
    input  logic       sd_clk_i        ,
    output logic [7:0] leds_o          ,
    input  logic [7:0] dip_switches_i
);

    // ---------------
    // 1. PLIC
    // ---------------
    logic [ariane_soc::NumSources-1:0] irq_sources;

    // Unused interrupt sources
    assign irq_sources[ariane_soc::NumSources-1:8] = '0;

    REG_BUS #(
        .ADDR_WIDTH ( 32 ),
        .DATA_WIDTH ( 32 )
    ) reg_bus (clk_i);

    logic         plic_penable;
    logic         plic_pwrite;
    logic [31:0]  plic_paddr;
    logic         plic_psel;
    logic [31:0]  plic_pwdata;
    logic [31:0]  plic_prdata;
    logic         plic_pready;
    logic         plic_pslverr;

    axi2apb_64_32 #(
        .AXI4_ADDRESS_WIDTH ( AxiAddrWidth  ),
        .AXI4_RDATA_WIDTH   ( AxiDataWidth  ),
        .AXI4_WDATA_WIDTH   ( AxiDataWidth  ),
        .AXI4_ID_WIDTH      ( AxiIdWidth    ),
        .AXI4_USER_WIDTH    ( AxiUserWidth  ),
        .BUFF_DEPTH_SLAVE   ( 2             ),
        .APB_ADDR_WIDTH     ( 32            )
    ) i_axi2apb_64_32_plic (
        .ACLK      ( clk_i          ),
        .ARESETn   ( rst_ni         ),
        .test_en_i ( 1'b0           ),
        .AWID_i    ( plic.aw_id     ),
        .AWADDR_i  ( plic.aw_addr   ),
        .AWLEN_i   ( plic.aw_len    ),
        .AWSIZE_i  ( plic.aw_size   ),
        .AWBURST_i ( plic.aw_burst  ),
        .AWLOCK_i  ( plic.aw_lock   ),
        .AWCACHE_i ( plic.aw_cache  ),
        .AWPROT_i  ( plic.aw_prot   ),
        .AWREGION_i( plic.aw_region ),
        .AWUSER_i  ( plic.aw_user   ),
        .AWQOS_i   ( plic.aw_qos    ),
        .AWVALID_i ( plic.aw_valid  ),
        .AWREADY_o ( plic.aw_ready  ),
        .WDATA_i   ( plic.w_data    ),
        .WSTRB_i   ( plic.w_strb    ),
        .WLAST_i   ( plic.w_last    ),
        .WUSER_i   ( plic.w_user    ),
        .WVALID_i  ( plic.w_valid   ),
        .WREADY_o  ( plic.w_ready   ),
        .BID_o     ( plic.b_id      ),
        .BRESP_o   ( plic.b_resp    ),
        .BVALID_o  ( plic.b_valid   ),
        .BUSER_o   ( plic.b_user    ),
        .BREADY_i  ( plic.b_ready   ),
        .ARID_i    ( plic.ar_id     ),
        .ARADDR_i  ( plic.ar_addr   ),
        .ARLEN_i   ( plic.ar_len    ),
        .ARSIZE_i  ( plic.ar_size   ),
        .ARBURST_i ( plic.ar_burst  ),
        .ARLOCK_i  ( plic.ar_lock   ),
        .ARCACHE_i ( plic.ar_cache  ),
        .ARPROT_i  ( plic.ar_prot   ),
        .ARREGION_i( plic.ar_region ),
        .ARUSER_i  ( plic.ar_user   ),
        .ARQOS_i   ( plic.ar_qos    ),
        .ARVALID_i ( plic.ar_valid  ),
        .ARREADY_o ( plic.ar_ready  ),
        .RID_o     ( plic.r_id      ),
        .RDATA_o   ( plic.r_data    ),
        .RRESP_o   ( plic.r_resp    ),
        .RLAST_o   ( plic.r_last    ),
        .RUSER_o   ( plic.r_user    ),
        .RVALID_o  ( plic.r_valid   ),
        .RREADY_i  ( plic.r_ready   ),
        .PENABLE   ( plic_penable   ),
        .PWRITE    ( plic_pwrite    ),
        .PADDR     ( plic_paddr     ),
        .PSEL      ( plic_psel      ),
        .PWDATA    ( plic_pwdata    ),
        .PRDATA    ( plic_prdata    ),
        .PREADY    ( plic_pready    ),
        .PSLVERR   ( plic_pslverr   )
    );

    apb_to_reg i_apb_to_reg (
        .clk_i     ( clk_i        ),
        .rst_ni    ( rst_ni       ),
        .penable_i ( plic_penable ),
        .pwrite_i  ( plic_pwrite  ),
        .paddr_i   ( plic_paddr   ),
        .psel_i    ( plic_psel    ),
        .pwdata_i  ( plic_pwdata  ),
        .prdata_o  ( plic_prdata  ),
        .pready_o  ( plic_pready  ),
        .pslverr_o ( plic_pslverr ),
        .reg_o     ( reg_bus      )
    );

    // define reg type according to REG_BUS above
    `REG_BUS_TYPEDEF_ALL(plic, logic[31:0], logic[31:0], logic[3:0])
    plic_req_t plic_req;
    plic_rsp_t plic_rsp;

    // assign REG_BUS.out to (req_t, rsp_t) pair
    `REG_BUS_ASSIGN_TO_REQ(plic_req, reg_bus)
    `REG_BUS_ASSIGN_FROM_RSP(reg_bus, plic_rsp)

    plic_top #(
      .N_SOURCE    ( ariane_soc::NumSources  ),
      .N_TARGET    ( ariane_soc::NumTargets  ),
      .MAX_PRIO    ( ariane_soc::MaxPriority ),
      .reg_req_t   ( plic_req_t              ),
      .reg_rsp_t   ( plic_rsp_t              )
    ) i_plic (
      .clk_i,
      .rst_ni,
      .req_i         ( plic_req    ),
      .resp_o        ( plic_rsp    ),
      .le_i          ( '0          ), // 0:level 1:edge
      .irq_sources_i ( irq_sources ),
      .eip_targets_o ( irq_o       )
    );

    // ---------------
    // 2. UART
    // ---------------
    logic         uart_penable;
    logic         uart_pwrite;
    logic [31:0]  uart_paddr;
    logic         uart_psel;
    logic [31:0]  uart_pwdata;
    logic [31:0]  uart_prdata;
    logic         uart_pready;
    logic         uart_pslverr;

    axi2apb_64_32 #(
        .AXI4_ADDRESS_WIDTH ( AxiAddrWidth ),
        .AXI4_RDATA_WIDTH   ( AxiDataWidth ),
        .AXI4_WDATA_WIDTH   ( AxiDataWidth ),
        .AXI4_ID_WIDTH      ( AxiIdWidth   ),
        .AXI4_USER_WIDTH    ( AxiUserWidth ),
        .BUFF_DEPTH_SLAVE   ( 2            ),
        .APB_ADDR_WIDTH     ( 32           )
    ) i_axi2apb_64_32_uart (
        .ACLK      ( clk_i          ),
        .ARESETn   ( rst_ni         ),
        .test_en_i ( 1'b0           ),
        .AWID_i    ( uart.aw_id     ),
        .AWADDR_i  ( uart.aw_addr   ),
        .AWLEN_i   ( uart.aw_len    ),
        .AWSIZE_i  ( uart.aw_size   ),
        .AWBURST_i ( uart.aw_burst  ),
        .AWLOCK_i  ( uart.aw_lock   ),
        .AWCACHE_i ( uart.aw_cache  ),
        .AWPROT_i  ( uart.aw_prot   ),
        .AWREGION_i( uart.aw_region ),
        .AWUSER_i  ( uart.aw_user   ),
        .AWQOS_i   ( uart.aw_qos    ),
        .AWVALID_i ( uart.aw_valid  ),
        .AWREADY_o ( uart.aw_ready  ),
        .WDATA_i   ( uart.w_data    ),
        .WSTRB_i   ( uart.w_strb    ),
        .WLAST_i   ( uart.w_last    ),
        .WUSER_i   ( uart.w_user    ),
        .WVALID_i  ( uart.w_valid   ),
        .WREADY_o  ( uart.w_ready   ),
        .BID_o     ( uart.b_id      ),
        .BRESP_o   ( uart.b_resp    ),
        .BVALID_o  ( uart.b_valid   ),
        .BUSER_o   ( uart.b_user    ),
        .BREADY_i  ( uart.b_ready   ),
        .ARID_i    ( uart.ar_id     ),
        .ARADDR_i  ( uart.ar_addr   ),
        .ARLEN_i   ( uart.ar_len    ),
        .ARSIZE_i  ( uart.ar_size   ),
        .ARBURST_i ( uart.ar_burst  ),
        .ARLOCK_i  ( uart.ar_lock   ),
        .ARCACHE_i ( uart.ar_cache  ),
        .ARPROT_i  ( uart.ar_prot   ),
        .ARREGION_i( uart.ar_region ),
        .ARUSER_i  ( uart.ar_user   ),
        .ARQOS_i   ( uart.ar_qos    ),
        .ARVALID_i ( uart.ar_valid  ),
        .ARREADY_o ( uart.ar_ready  ),
        .RID_o     ( uart.r_id      ),
        .RDATA_o   ( uart.r_data    ),
        .RRESP_o   ( uart.r_resp    ),
        .RLAST_o   ( uart.r_last    ),
        .RUSER_o   ( uart.r_user    ),
        .RVALID_o  ( uart.r_valid   ),
        .RREADY_i  ( uart.r_ready   ),
        .PENABLE   ( uart_penable   ),
        .PWRITE    ( uart_pwrite    ),
        .PADDR     ( uart_paddr     ),
        .PSEL      ( uart_psel      ),
        .PWDATA    ( uart_pwdata    ),
        .PRDATA    ( uart_prdata    ),
        .PREADY    ( uart_pready    ),
        .PSLVERR   ( uart_pslverr   )
    );

    if (InclUART) begin : gen_uart
        apb_uart i_apb_uart (
            .CLK     ( clk_i           ),
            .RSTN    ( rst_ni          ),
            .PSEL    ( uart_psel       ),
            .PENABLE ( uart_penable    ),
            .PWRITE  ( uart_pwrite     ),
            .PADDR   ( uart_paddr[4:2] ),
            .PWDATA  ( uart_pwdata     ),
            .PRDATA  ( uart_prdata     ),
            .PREADY  ( uart_pready     ),
            .PSLVERR ( uart_pslverr    ),
            .INT     ( irq_sources[0]  ),
            .OUT1N   (                 ), // keep open
            .OUT2N   (                 ), // keep open
            .RTSN    (                 ), // no flow control
            .DTRN    (                 ), // no flow control
            .CTSN    ( 1'b0            ),
            .DSRN    ( 1'b0            ),
            .DCDN    ( 1'b0            ),
            .RIN     ( 1'b0            ),
            .SIN     ( rx_i            ),
            .SOUT    ( tx_o            )
        );
    end else begin
        /* pragma translate_off */
        `ifndef VERILATOR
        mock_uart i_mock_uart (
            .clk_i     ( clk_i        ),
            .rst_ni    ( rst_ni       ),
            .penable_i ( uart_penable ),
            .pwrite_i  ( uart_pwrite  ),
            .paddr_i   ( uart_paddr   ),
            .psel_i    ( uart_psel    ),
            .pwdata_i  ( uart_pwdata  ),
            .prdata_o  ( uart_prdata  ),
            .pready_o  ( uart_pready  ),
            .pslverr_o ( uart_pslverr )
        );
        `endif
        /* pragma translate_on */
    end

    // ---------------
    // 3. SPI
    // ---------------
    assign spi.b_user = 1'b0;
    assign spi.r_user = 1'b0;

    if (InclSPI) begin : gen_spi
        logic [31:0] s_axi_spi_awaddr;
        logic [7:0]  s_axi_spi_awlen;
        logic [2:0]  s_axi_spi_awsize;
        logic [1:0]  s_axi_spi_awburst;
        logic [0:0]  s_axi_spi_awlock;
        logic [3:0]  s_axi_spi_awcache;
        logic [2:0]  s_axi_spi_awprot;
        logic [3:0]  s_axi_spi_awregion;
        logic [3:0]  s_axi_spi_awqos;
        logic        s_axi_spi_awvalid;
        logic        s_axi_spi_awready;
        logic [31:0] s_axi_spi_wdata;
        logic [3:0]  s_axi_spi_wstrb;
        logic        s_axi_spi_wlast;
        logic        s_axi_spi_wvalid;
        logic        s_axi_spi_wready;
        logic [1:0]  s_axi_spi_bresp;
        logic        s_axi_spi_bvalid;
        logic        s_axi_spi_bready;
        logic [31:0] s_axi_spi_araddr;
        logic [7:0]  s_axi_spi_arlen;
        logic [2:0]  s_axi_spi_arsize;
        logic [1:0]  s_axi_spi_arburst;
        logic [0:0]  s_axi_spi_arlock;
        logic [3:0]  s_axi_spi_arcache;
        logic [2:0]  s_axi_spi_arprot;
        logic [3:0]  s_axi_spi_arregion;
        logic [3:0]  s_axi_spi_arqos;
        logic        s_axi_spi_arvalid;
        logic        s_axi_spi_arready;
        logic [31:0] s_axi_spi_rdata;
        logic [1:0]  s_axi_spi_rresp;
        logic        s_axi_spi_rlast;
        logic        s_axi_spi_rvalid;
        logic        s_axi_spi_rready;

        xlnx_axi_dwidth_converter i_xlnx_axi_dwidth_converter_spi (
            .s_axi_aclk     ( clk_i              ),
            .s_axi_aresetn  ( rst_ni             ),

            .s_axi_awid     ( spi.aw_id          ),
            .s_axi_awaddr   ( spi.aw_addr[31:0]  ),
            .s_axi_awlen    ( spi.aw_len         ),
            .s_axi_awsize   ( spi.aw_size        ),
            .s_axi_awburst  ( spi.aw_burst       ),
            .s_axi_awlock   ( spi.aw_lock        ),
            .s_axi_awcache  ( spi.aw_cache       ),
            .s_axi_awprot   ( spi.aw_prot        ),
            .s_axi_awregion ( spi.aw_region      ),
            .s_axi_awqos    ( spi.aw_qos         ),
            .s_axi_awvalid  ( spi.aw_valid       ),
            .s_axi_awready  ( spi.aw_ready       ),
            .s_axi_wdata    ( spi.w_data         ),
            .s_axi_wstrb    ( spi.w_strb         ),
            .s_axi_wlast    ( spi.w_last         ),
            .s_axi_wvalid   ( spi.w_valid        ),
            .s_axi_wready   ( spi.w_ready        ),
            .s_axi_bid      ( spi.b_id           ),
            .s_axi_bresp    ( spi.b_resp         ),
            .s_axi_bvalid   ( spi.b_valid        ),
            .s_axi_bready   ( spi.b_ready        ),
            .s_axi_arid     ( spi.ar_id          ),
            .s_axi_araddr   ( spi.ar_addr[31:0]  ),
            .s_axi_arlen    ( spi.ar_len         ),
            .s_axi_arsize   ( spi.ar_size        ),
            .s_axi_arburst  ( spi.ar_burst       ),
            .s_axi_arlock   ( spi.ar_lock        ),
            .s_axi_arcache  ( spi.ar_cache       ),
            .s_axi_arprot   ( spi.ar_prot        ),
            .s_axi_arregion ( spi.ar_region      ),
            .s_axi_arqos    ( spi.ar_qos         ),
            .s_axi_arvalid  ( spi.ar_valid       ),
            .s_axi_arready  ( spi.ar_ready       ),
            .s_axi_rid      ( spi.r_id           ),
            .s_axi_rdata    ( spi.r_data         ),
            .s_axi_rresp    ( spi.r_resp         ),
            .s_axi_rlast    ( spi.r_last         ),
            .s_axi_rvalid   ( spi.r_valid        ),
            .s_axi_rready   ( spi.r_ready        ),

            .m_axi_awaddr   ( s_axi_spi_awaddr   ),
            .m_axi_awlen    ( s_axi_spi_awlen    ),
            .m_axi_awsize   ( s_axi_spi_awsize   ),
            .m_axi_awburst  ( s_axi_spi_awburst  ),
            .m_axi_awlock   ( s_axi_spi_awlock   ),
            .m_axi_awcache  ( s_axi_spi_awcache  ),
            .m_axi_awprot   ( s_axi_spi_awprot   ),
            .m_axi_awregion ( s_axi_spi_awregion ),
            .m_axi_awqos    ( s_axi_spi_awqos    ),
            .m_axi_awvalid  ( s_axi_spi_awvalid  ),
            .m_axi_awready  ( s_axi_spi_awready  ),
            .m_axi_wdata    ( s_axi_spi_wdata    ),
            .m_axi_wstrb    ( s_axi_spi_wstrb    ),
            .m_axi_wlast    ( s_axi_spi_wlast    ),
            .m_axi_wvalid   ( s_axi_spi_wvalid   ),
            .m_axi_wready   ( s_axi_spi_wready   ),
            .m_axi_bresp    ( s_axi_spi_bresp    ),
            .m_axi_bvalid   ( s_axi_spi_bvalid   ),
            .m_axi_bready   ( s_axi_spi_bready   ),
            .m_axi_araddr   ( s_axi_spi_araddr   ),
            .m_axi_arlen    ( s_axi_spi_arlen    ),
            .m_axi_arsize   ( s_axi_spi_arsize   ),
            .m_axi_arburst  ( s_axi_spi_arburst  ),
            .m_axi_arlock   ( s_axi_spi_arlock   ),
            .m_axi_arcache  ( s_axi_spi_arcache  ),
            .m_axi_arprot   ( s_axi_spi_arprot   ),
            .m_axi_arregion ( s_axi_spi_arregion ),
            .m_axi_arqos    ( s_axi_spi_arqos    ),
            .m_axi_arvalid  ( s_axi_spi_arvalid  ),
            .m_axi_arready  ( s_axi_spi_arready  ),
            .m_axi_rdata    ( s_axi_spi_rdata    ),
            .m_axi_rresp    ( s_axi_spi_rresp    ),
            .m_axi_rlast    ( s_axi_spi_rlast    ),
            .m_axi_rvalid   ( s_axi_spi_rvalid   ),
            .m_axi_rready   ( s_axi_spi_rready   )
        );

        xlnx_axi_quad_spi i_xlnx_axi_quad_spi (
            .ext_spi_clk    ( clk_i                  ),
            .s_axi4_aclk    ( clk_i                  ),
            .s_axi4_aresetn ( rst_ni                 ),
            .s_axi4_awaddr  ( s_axi_spi_awaddr[23:0] ),
            .s_axi4_awlen   ( s_axi_spi_awlen        ),
            .s_axi4_awsize  ( s_axi_spi_awsize       ),
            .s_axi4_awburst ( s_axi_spi_awburst      ),
            .s_axi4_awlock  ( s_axi_spi_awlock       ),
            .s_axi4_awcache ( s_axi_spi_awcache      ),
            .s_axi4_awprot  ( s_axi_spi_awprot       ),
            .s_axi4_awvalid ( s_axi_spi_awvalid      ),
            .s_axi4_awready ( s_axi_spi_awready      ),
            .s_axi4_wdata   ( s_axi_spi_wdata        ),
            .s_axi4_wstrb   ( s_axi_spi_wstrb        ),
            .s_axi4_wlast   ( s_axi_spi_wlast        ),
            .s_axi4_wvalid  ( s_axi_spi_wvalid       ),
            .s_axi4_wready  ( s_axi_spi_wready       ),
            .s_axi4_bresp   ( s_axi_spi_bresp        ),
            .s_axi4_bvalid  ( s_axi_spi_bvalid       ),
            .s_axi4_bready  ( s_axi_spi_bready       ),
            .s_axi4_araddr  ( s_axi_spi_araddr[23:0] ),
            .s_axi4_arlen   ( s_axi_spi_arlen        ),
            .s_axi4_arsize  ( s_axi_spi_arsize       ),
            .s_axi4_arburst ( s_axi_spi_arburst      ),
            .s_axi4_arlock  ( s_axi_spi_arlock       ),
            .s_axi4_arcache ( s_axi_spi_arcache      ),
            .s_axi4_arprot  ( s_axi_spi_arprot       ),
            .s_axi4_arvalid ( s_axi_spi_arvalid      ),
            .s_axi4_arready ( s_axi_spi_arready      ),
            .s_axi4_rdata   ( s_axi_spi_rdata        ),
            .s_axi4_rresp   ( s_axi_spi_rresp        ),
            .s_axi4_rlast   ( s_axi_spi_rlast        ),
            .s_axi4_rvalid  ( s_axi_spi_rvalid       ),
            .s_axi4_rready  ( s_axi_spi_rready       ),
            .io0_i          ( '0                     ),
            .io0_o          ( spi_mosi               ),
            .io0_t          (                        ),
            .io1_i          ( spi_miso               ),
            .io1_o          (                        ),
            .io1_t          (                        ),
            .ss_i           ( '0                     ),
            .ss_o           ( spi_ss                 ),
            .ss_t           (                        ),
            .sck_o          ( spi_clk_o              ),
            .sck_i          ( '0                     ),
            .sck_t          (                        ),
            .ip2intc_irpt   ( irq_sources[1]         )
        );
    end else begin
        assign spi_clk_o = 1'b0;
        assign spi_mosi = 1'b0;
        assign spi_ss = 1'b0;

        // assign irq_sources [1] = 1'b0;
        assign spi.aw_ready = 1'b1;
        assign spi.ar_ready = 1'b1;
        assign spi.w_ready = 1'b1;

        assign spi.b_valid = spi.aw_valid;
        assign spi.b_id = spi.aw_id;
        assign spi.b_resp = axi_pkg::RESP_SLVERR;
        assign spi.b_user = '0;

        assign spi.r_valid = spi.ar_valid;
        assign spi.r_resp = axi_pkg::RESP_SLVERR;
        assign spi.r_data = 'hdeadbeef;
        assign spi.r_last = 1'b1;
    end


    // ---------------
    // 4. Ethernet
    // ---------------

    if (InclXilinxEthernet || InclLowriscEthernet) begin : gen_ethernet_common
        // Code common to both Ethernet MACs.

        logic eth_mdio_i, eth_mdio_o, eth_mdio_oe;

        IOBUF #(
           .DRIVE(12), // Specify the output drive strength
           .IBUF_LOW_PWR("TRUE"),  // Low Power - "TRUE", High Performance = "FALSE"
           .IOSTANDARD("DEFAULT"), // Specify the I/O standard
           .SLEW("SLOW") // Specify the output slew rate
        ) IOBUF_inst (
           .O(eth_mdio_i),     // Buffer output
           .IO(eth_mdio),   // Buffer inout port (connect directly to top-level port)
           .I(eth_mdio_o),     // Buffer input
           .T(eth_mdio_oe)      // 3-state enable input, high=input, low=output
        );

    end else begin
        // Tie off signals with no ethernet
        assign irq_sources [2] = 1'b0;
        assign ethernet_data.aw_ready = 1'b1;
        assign ethernet_data.ar_ready = 1'b1;
        assign ethernet_data.w_ready = 1'b1;

        assign ethernet_data.b_valid = ethernet_data.aw_valid;
        assign ethernet_data.b_id = ethernet_data.aw_id;
        assign ethernet_data.b_resp = axi_pkg::RESP_SLVERR;
        assign ethernet_data.b_user = '0;

        assign ethernet_data.r_valid = ethernet_data.ar_valid;
        assign ethernet_data.r_resp = axi_pkg::RESP_SLVERR;
        assign ethernet_data.r_data = 'hdeadbeef;
        assign ethernet_data.r_last = 1'b1;
    end

    if (InclXilinxEthernet) begin : gen_axi_ethernet
        // Convert the incoming ethernet FIFO master down to 32bits
        logic [31:0] s_axi_ethernet_data_awaddr;
        logic [7:0]  s_axi_ethernet_data_awlen;
        logic [2:0]  s_axi_ethernet_data_awsize;
        logic [1:0]  s_axi_ethernet_data_awburst;
        logic [0:0]  s_axi_ethernet_data_awlock;
        logic [3:0]  s_axi_ethernet_data_awcache;
        logic [2:0]  s_axi_ethernet_data_awprot;
        logic [3:0]  s_axi_ethernet_data_awregion;
        logic [3:0]  s_axi_ethernet_data_awqos;
        logic        s_axi_ethernet_data_awvalid;
        logic        s_axi_ethernet_data_awready;
        logic [31:0] s_axi_ethernet_data_wdata;
        logic [3:0]  s_axi_ethernet_data_wstrb;
        logic        s_axi_ethernet_data_wlast;
        logic        s_axi_ethernet_data_wvalid;
        logic        s_axi_ethernet_data_wready;
        logic [1:0]  s_axi_ethernet_data_bresp;
        logic        s_axi_ethernet_data_bvalid;
        logic        s_axi_ethernet_data_bready;
        logic [31:0] s_axi_ethernet_data_araddr;
        logic [7:0]  s_axi_ethernet_data_arlen;
        logic [2:0]  s_axi_ethernet_data_arsize;
        logic [1:0]  s_axi_ethernet_data_arburst;
        logic [0:0]  s_axi_ethernet_data_arlock;
        logic [3:0]  s_axi_ethernet_data_arcache;
        logic [2:0]  s_axi_ethernet_data_arprot;
        logic [3:0]  s_axi_ethernet_data_arregion;
        logic [3:0]  s_axi_ethernet_data_arqos;
        logic        s_axi_ethernet_data_arvalid;
        logic        s_axi_ethernet_data_arready;
        logic [31:0] s_axi_ethernet_data_rdata;
        logic [1:0]  s_axi_ethernet_data_rresp;
        logic        s_axi_ethernet_data_rlast;
        logic        s_axi_ethernet_data_rvalid;
        logic        s_axi_ethernet_data_rready;

        xlnx_axi_dwidth_converter i_xlnx_axi_dwidth_converter_ethernet_data (
            .s_axi_aclk     ( clk_i                        ),
            .s_axi_aresetn  ( rst_ni                       ),

            .s_axi_awid     ( ethernet_data.aw_id          ),
            .s_axi_awaddr   ( ethernet_data.aw_addr[31:0]  ),
            .s_axi_awlen    ( ethernet_data.aw_len         ),
            .s_axi_awsize   ( ethernet_data.aw_size        ),
            .s_axi_awburst  ( ethernet_data.aw_burst       ),
            .s_axi_awlock   ( ethernet_data.aw_lock        ),
            .s_axi_awcache  ( ethernet_data.aw_cache       ),
            .s_axi_awprot   ( ethernet_data.aw_prot        ),
            .s_axi_awregion ( ethernet_data.aw_region      ),
            .s_axi_awqos    ( ethernet_data.aw_qos         ),
            .s_axi_awvalid  ( ethernet_data.aw_valid       ),
            .s_axi_awready  ( ethernet_data.aw_ready       ),
            .s_axi_wdata    ( ethernet_data.w_data         ),
            .s_axi_wstrb    ( ethernet_data.w_strb         ),
            .s_axi_wlast    ( ethernet_data.w_last         ),
            .s_axi_wvalid   ( ethernet_data.w_valid        ),
            .s_axi_wready   ( ethernet_data.w_ready        ),
            .s_axi_bid      ( ethernet_data.b_id           ),
            .s_axi_bresp    ( ethernet_data.b_resp         ),
            .s_axi_bvalid   ( ethernet_data.b_valid        ),
            .s_axi_bready   ( ethernet_data.b_ready        ),
            .s_axi_arid     ( ethernet_data.ar_id          ),
            .s_axi_araddr   ( ethernet_data.ar_addr[31:0]  ),
            .s_axi_arlen    ( ethernet_data.ar_len         ),
            .s_axi_arsize   ( ethernet_data.ar_size        ),
            .s_axi_arburst  ( ethernet_data.ar_burst       ),
            .s_axi_arlock   ( ethernet_data.ar_lock        ),
            .s_axi_arcache  ( ethernet_data.ar_cache       ),
            .s_axi_arprot   ( ethernet_data.ar_prot        ),
            .s_axi_arregion ( ethernet_data.ar_region      ),
            .s_axi_arqos    ( ethernet_data.ar_qos         ),
            .s_axi_arvalid  ( ethernet_data.ar_valid       ),
            .s_axi_arready  ( ethernet_data.ar_ready       ),
            .s_axi_rid      ( ethernet_data.r_id           ),
            .s_axi_rdata    ( ethernet_data.r_data         ),
            .s_axi_rresp    ( ethernet_data.r_resp         ),
            .s_axi_rlast    ( ethernet_data.r_last         ),
            .s_axi_rvalid   ( ethernet_data.r_valid        ),
            .s_axi_rready   ( ethernet_data.r_ready        ),

            .m_axi_awaddr   ( s_axi_ethernet_data_awaddr   ),
            .m_axi_awlen    ( s_axi_ethernet_data_awlen    ),
            .m_axi_awsize   ( s_axi_ethernet_data_awsize   ),
            .m_axi_awburst  ( s_axi_ethernet_data_awburst  ),
            .m_axi_awlock   ( s_axi_ethernet_data_awlock   ),
            .m_axi_awcache  ( s_axi_ethernet_data_awcache  ),
            .m_axi_awprot   ( s_axi_ethernet_data_awprot   ),
            .m_axi_awregion ( s_axi_ethernet_data_awregion ),
            .m_axi_awqos    ( s_axi_ethernet_data_awqos    ),
            .m_axi_awvalid  ( s_axi_ethernet_data_awvalid  ),
            .m_axi_awready  ( s_axi_ethernet_data_awready  ),
            .m_axi_wdata    ( s_axi_ethernet_data_wdata    ),
            .m_axi_wstrb    ( s_axi_ethernet_data_wstrb    ),
            .m_axi_wlast    ( s_axi_ethernet_data_wlast    ),
            .m_axi_wvalid   ( s_axi_ethernet_data_wvalid   ),
            .m_axi_wready   ( s_axi_ethernet_data_wready   ),
            .m_axi_bresp    ( s_axi_ethernet_data_bresp    ),
            .m_axi_bvalid   ( s_axi_ethernet_data_bvalid   ),
            .m_axi_bready   ( s_axi_ethernet_data_bready   ),
            .m_axi_araddr   ( s_axi_ethernet_data_araddr   ),
            .m_axi_arlen    ( s_axi_ethernet_data_arlen    ),
            .m_axi_arsize   ( s_axi_ethernet_data_arsize   ),
            .m_axi_arburst  ( s_axi_ethernet_data_arburst  ),
            .m_axi_arlock   ( s_axi_ethernet_data_arlock   ),
            .m_axi_arcache  ( s_axi_ethernet_data_arcache  ),
            .m_axi_arprot   ( s_axi_ethernet_data_arprot   ),
            .m_axi_arregion ( s_axi_ethernet_data_arregion ),
            .m_axi_arqos    ( s_axi_ethernet_data_arqos    ),
            .m_axi_arvalid  ( s_axi_ethernet_data_arvalid  ),
            .m_axi_arready  ( s_axi_ethernet_data_arready  ),
            .m_axi_rdata    ( s_axi_ethernet_data_rdata    ),
            .m_axi_rresp    ( s_axi_ethernet_data_rresp    ),
            .m_axi_rlast    ( s_axi_ethernet_data_rlast    ),
            .m_axi_rvalid   ( s_axi_ethernet_data_rvalid   ),
            .m_axi_rready   ( s_axi_ethernet_data_rready   )
        );

        // Convert the full AXI ethernet FIFO master into AXI lite
        logic [31:0] s_axi_lite_ethernet_data_awaddr;
        logic        s_axi_lite_ethernet_data_awvalid;
        logic        s_axi_lite_ethernet_data_awready;
        logic [31:0] s_axi_lite_ethernet_data_wdata;
        logic [3:0]  s_axi_lite_ethernet_data_wstrb;
        logic        s_axi_lite_ethernet_data_wvalid;
        logic        s_axi_lite_ethernet_data_wready;
        logic [1:0]  s_axi_lite_ethernet_data_bresp;
        logic        s_axi_lite_ethernet_data_bvalid;
        logic        s_axi_lite_ethernet_data_bready;
        logic [31:0] s_axi_lite_ethernet_data_araddr;
        logic        s_axi_lite_ethernet_data_arvalid;
        logic        s_axi_lite_ethernet_data_arready;
        logic [31:0] s_axi_lite_ethernet_data_rdata;
        logic [1:0]  s_axi_lite_ethernet_data_rresp;
        logic        s_axi_lite_ethernet_data_rvalid;
        logic        s_axi_lite_ethernet_data_rready;

        xlnx_axi_lite_converter i_xlnx_axi_lite_converter_ethernet_data (
            .aclk           ( clk_i                            ),
            .aresetn        ( rst_ni                           ),

            .s_axi_awaddr   ( s_axi_ethernet_data_awaddr       ),
            .s_axi_awlen    ( s_axi_ethernet_data_awlen        ),
            .s_axi_awsize   ( s_axi_ethernet_data_awsize       ),
            .s_axi_awburst  ( s_axi_ethernet_data_awburst      ),
            .s_axi_awlock   ( s_axi_ethernet_data_awlock       ),
            .s_axi_awcache  ( s_axi_ethernet_data_awcache      ),
            .s_axi_awprot   ( s_axi_ethernet_data_awprot       ),
            .s_axi_awregion ( s_axi_ethernet_data_awregion     ),
            .s_axi_awqos    ( s_axi_ethernet_data_awqos        ),
            .s_axi_awvalid  ( s_axi_ethernet_data_awvalid      ),
            .s_axi_awready  ( s_axi_ethernet_data_awready      ),
            .s_axi_wdata    ( s_axi_ethernet_data_wdata        ),
            .s_axi_wstrb    ( s_axi_ethernet_data_wstrb        ),
            .s_axi_wlast    ( s_axi_ethernet_data_wlast        ),
            .s_axi_wvalid   ( s_axi_ethernet_data_wvalid       ),
            .s_axi_wready   ( s_axi_ethernet_data_wready       ),
            .s_axi_bresp    ( s_axi_ethernet_data_bresp        ),
            .s_axi_bvalid   ( s_axi_ethernet_data_bvalid       ),
            .s_axi_bready   ( s_axi_ethernet_data_bready       ),
            .s_axi_araddr   ( s_axi_ethernet_data_araddr       ),
            .s_axi_arlen    ( s_axi_ethernet_data_arlen        ),
            .s_axi_arsize   ( s_axi_ethernet_data_arsize       ),
            .s_axi_arburst  ( s_axi_ethernet_data_arburst      ),
            .s_axi_arlock   ( s_axi_ethernet_data_arlock       ),
            .s_axi_arcache  ( s_axi_ethernet_data_arcache      ),
            .s_axi_arprot   ( s_axi_ethernet_data_arprot       ),
            .s_axi_arregion ( s_axi_ethernet_data_arregion     ),
            .s_axi_arqos    ( s_axi_ethernet_data_arqos        ),
            .s_axi_arvalid  ( s_axi_ethernet_data_arvalid      ),
            .s_axi_arready  ( s_axi_ethernet_data_arready      ),
            .s_axi_rdata    ( s_axi_ethernet_data_rdata        ),
            .s_axi_rresp    ( s_axi_ethernet_data_rresp        ),
            .s_axi_rlast    ( s_axi_ethernet_data_rlast        ),
            .s_axi_rvalid   ( s_axi_ethernet_data_rvalid       ),
            .s_axi_rready   ( s_axi_ethernet_data_rready       ),

            .m_axi_awaddr   ( s_axi_lite_ethernet_data_awaddr  ),
            .m_axi_awprot   ( /* NC */                         ),
            .m_axi_awvalid  ( s_axi_lite_ethernet_data_awvalid ),
            .m_axi_awready  ( s_axi_lite_ethernet_data_awready ),
            .m_axi_wdata    ( s_axi_lite_ethernet_data_wdata   ),
            .m_axi_wstrb    ( s_axi_lite_ethernet_data_wstrb   ),
            .m_axi_wvalid   ( s_axi_lite_ethernet_data_wvalid  ),
            .m_axi_wready   ( s_axi_lite_ethernet_data_wready  ),
            .m_axi_bresp    ( s_axi_lite_ethernet_data_bresp   ),
            .m_axi_bvalid   ( s_axi_lite_ethernet_data_bvalid  ),
            .m_axi_bready   ( s_axi_lite_ethernet_data_bready  ),
            .m_axi_araddr   ( s_axi_lite_ethernet_data_araddr  ),
            .m_axi_arprot   ( /* NC */                         ),
            .m_axi_arvalid  ( s_axi_lite_ethernet_data_arvalid ),
            .m_axi_arready  ( s_axi_lite_ethernet_data_arready ),
            .m_axi_rdata    ( s_axi_lite_ethernet_data_rdata   ),
            .m_axi_rresp    ( s_axi_lite_ethernet_data_rresp   ),
            .m_axi_rvalid   ( s_axi_lite_ethernet_data_rvalid  ),
            .m_axi_rready   ( s_axi_lite_ethernet_data_rready  )
        );

        logic        mm2s_prmry_reset_out_n;
        logic        fifo_axi_str_txd_tvalid;
        logic        fifo_axi_str_txd_tready;
        logic        fifo_axi_str_txd_tlast;
        logic [3:0]  fifo_axi_str_txd_tkeep;
        logic [31:0] fifo_axi_str_txd_tdata;
        logic        fifo_mm2s_cntrl_reset_out_n;
        logic        fifo_axi_str_txc_tvalid;
        logic        fifo_axi_str_txc_tready;
        logic        fifo_axi_str_txc_tlast;
        logic [3:0]  fifo_axi_str_txc_tkeep;
        logic [31:0] fifo_axi_str_txc_tdata;
        logic        fifo_s2mm_prmry_reset_out_n;
        logic        fifo_axi_str_rxd_tvalid;
        logic        fifo_axi_str_rxd_tready;
        logic        fifo_axi_str_rxd_tlast;
        logic [3:0]  fifo_axi_str_rxd_tkeep;
        logic [31:0] fifo_axi_str_rxd_tdata;

        xlnx_axi_fifo (
            .interrupt              ( irq_sources[7]                   ),
            .s_axi_aclk             ( clk_i                            ),
            .s_axi_aresetn          ( rst_ni                           ),
            .s_axi_awaddr           ( s_axi_lite_ethernet_data_awaddr  ),
            .s_axi_awvalid          ( s_axi_lite_ethernet_data_awvalid ),
            .s_axi_awready          ( s_axi_lite_ethernet_data_awready ),
            .s_axi_wdata            ( s_axi_lite_ethernet_data_wdata   ),
            .s_axi_wstrb            ( s_axi_lite_ethernet_data_wstrb   ),
            .s_axi_wvalid           ( s_axi_lite_ethernet_data_wvalid  ),
            .s_axi_wready           ( s_axi_lite_ethernet_data_wready  ),
            .s_axi_bresp            ( s_axi_lite_ethernet_data_bresp   ),
            .s_axi_bvalid           ( s_axi_lite_ethernet_data_bvalid  ),
            .s_axi_bready           ( s_axi_lite_ethernet_data_bready  ),
            .s_axi_araddr           ( s_axi_lite_ethernet_data_araddr  ),
            .s_axi_arvalid          ( s_axi_lite_ethernet_data_arvalid ),
            .s_axi_arready          ( s_axi_lite_ethernet_data_arready ),
            .s_axi_rdata            ( s_axi_lite_ethernet_data_rdata   ),
            .s_axi_rresp            ( s_axi_lite_ethernet_data_rresp   ),
            .s_axi_rvalid           ( s_axi_lite_ethernet_data_rvalid  ),
            .s_axi_rready           ( s_axi_lite_ethernet_data_rready  ),
            .mm2s_prmry_reset_out_n ( fifo_mm2s_prmry_reset_out_n      ),
            .axi_str_txd_tvalid     ( fifo_axi_str_txd_tvalid          ),
            .axi_str_txd_tready     ( fifo_axi_str_txd_tready          ),
            .axi_str_txd_tlast      ( fifo_axi_str_txd_tlast           ),
            .axi_str_txd_tkeep      ( fifo_axi_str_txd_tkeep           ),
            .axi_str_txd_tdata      ( fifo_axi_str_txd_tdata           ),
            .mm2s_cntrl_reset_out_n ( fifo_mm2s_cntrl_reset_out_n      ),
            .axi_str_txc_tvalid     ( fifo_axi_str_txc_tvalid          ),
            .axi_str_txc_tready     ( fifo_axi_str_txc_tready          ),
            .axi_str_txc_tlast      ( fifo_axi_str_txc_tlast           ),
            .axi_str_txc_tkeep      ( fifo_axi_str_txc_tkeep           ),
            .axi_str_txc_tdata      ( fifo_axi_str_txc_tdata           ),
            .s2mm_prmry_reset_out_n ( fifo_s2mm_prmry_reset_out_n      ),
            .axi_str_rxd_tvalid     ( fifo_axi_str_rxd_tvalid          ),
            .axi_str_rxd_tready     ( fifo_axi_str_rxd_tready          ),
            .axi_str_rxd_tlast      ( fifo_axi_str_rxd_tlast           ),
            .axi_str_rxd_tkeep      ( fifo_axi_str_rxd_tkeep           ),
            .axi_str_rxd_tdata      ( fifo_axi_str_rxd_tdata           )
        );

        // Convert the incoming ethernet MAC master down to 32bits
        logic [31:0] s_axi_ethernet_mgmt_awaddr;
        logic [7:0]  s_axi_ethernet_mgmt_awlen;
        logic [2:0]  s_axi_ethernet_mgmt_awsize;
        logic [1:0]  s_axi_ethernet_mgmt_awburst;
        logic [0:0]  s_axi_ethernet_mgmt_awlock;
        logic [3:0]  s_axi_ethernet_mgmt_awcache;
        logic [2:0]  s_axi_ethernet_mgmt_awprot;
        logic [3:0]  s_axi_ethernet_mgmt_awregion;
        logic [3:0]  s_axi_ethernet_mgmt_awqos;
        logic        s_axi_ethernet_mgmt_awvalid;
        logic        s_axi_ethernet_mgmt_awready;
        logic [31:0] s_axi_ethernet_mgmt_wdata;
        logic [3:0]  s_axi_ethernet_mgmt_wstrb;
        logic        s_axi_ethernet_mgmt_wlast;
        logic        s_axi_ethernet_mgmt_wvalid;
        logic        s_axi_ethernet_mgmt_wready;
        logic [1:0]  s_axi_ethernet_mgmt_bresp;
        logic        s_axi_ethernet_mgmt_bvalid;
        logic        s_axi_ethernet_mgmt_bready;
        logic [31:0] s_axi_ethernet_mgmt_araddr;
        logic [7:0]  s_axi_ethernet_mgmt_arlen;
        logic [2:0]  s_axi_ethernet_mgmt_arsize;
        logic [1:0]  s_axi_ethernet_mgmt_arburst;
        logic [0:0]  s_axi_ethernet_mgmt_arlock;
        logic [3:0]  s_axi_ethernet_mgmt_arcache;
        logic [2:0]  s_axi_ethernet_mgmt_arprot;
        logic [3:0]  s_axi_ethernet_mgmt_arregion;
        logic [3:0]  s_axi_ethernet_mgmt_arqos;
        logic        s_axi_ethernet_mgmt_arvalid;
        logic        s_axi_ethernet_mgmt_arready;
        logic [31:0] s_axi_ethernet_mgmt_rdata;
        logic [1:0]  s_axi_ethernet_mgmt_rresp;
        logic        s_axi_ethernet_mgmt_rlast;
        logic        s_axi_ethernet_mgmt_rvalid;
        logic        s_axi_ethernet_mgmt_rready;

        xlnx_axi_dwidth_converter i_xlnx_axi_dwidth_converter_ethernet_mgmt (
            .s_axi_aclk     ( clk_i                        ),
            .s_axi_aresetn  ( rst_ni                       ),

            .s_axi_awid     ( ethernet_mgmt.aw_id          ),
            .s_axi_awaddr   ( ethernet_mgmt.aw_addr[31:0]  ),
            .s_axi_awlen    ( ethernet_mgmt.aw_len         ),
            .s_axi_awsize   ( ethernet_mgmt.aw_size        ),
            .s_axi_awburst  ( ethernet_mgmt.aw_burst       ),
            .s_axi_awlock   ( ethernet_mgmt.aw_lock        ),
            .s_axi_awcache  ( ethernet_mgmt.aw_cache       ),
            .s_axi_awprot   ( ethernet_mgmt.aw_prot        ),
            .s_axi_awregion ( ethernet_mgmt.aw_region      ),
            .s_axi_awqos    ( ethernet_mgmt.aw_qos         ),
            .s_axi_awvalid  ( ethernet_mgmt.aw_valid       ),
            .s_axi_awready  ( ethernet_mgmt.aw_ready       ),
            .s_axi_wdata    ( ethernet_mgmt.w_data         ),
            .s_axi_wstrb    ( ethernet_mgmt.w_strb         ),
            .s_axi_wlast    ( ethernet_mgmt.w_last         ),
            .s_axi_wvalid   ( ethernet_mgmt.w_valid        ),
            .s_axi_wready   ( ethernet_mgmt.w_ready        ),
            .s_axi_bid      ( ethernet_mgmt.b_id           ),
            .s_axi_bresp    ( ethernet_mgmt.b_resp         ),
            .s_axi_bvalid   ( ethernet_mgmt.b_valid        ),
            .s_axi_bready   ( ethernet_mgmt.b_ready        ),
            .s_axi_arid     ( ethernet_mgmt.ar_id          ),
            .s_axi_araddr   ( ethernet_mgmt.ar_addr[31:0]  ),
            .s_axi_arlen    ( ethernet_mgmt.ar_len         ),
            .s_axi_arsize   ( ethernet_mgmt.ar_size        ),
            .s_axi_arburst  ( ethernet_mgmt.ar_burst       ),
            .s_axi_arlock   ( ethernet_mgmt.ar_lock        ),
            .s_axi_arcache  ( ethernet_mgmt.ar_cache       ),
            .s_axi_arprot   ( ethernet_mgmt.ar_prot        ),
            .s_axi_arregion ( ethernet_mgmt.ar_region      ),
            .s_axi_arqos    ( ethernet_mgmt.ar_qos         ),
            .s_axi_arvalid  ( ethernet_mgmt.ar_valid       ),
            .s_axi_arready  ( ethernet_mgmt.ar_ready       ),
            .s_axi_rid      ( ethernet_mgmt.r_id           ),
            .s_axi_rdata    ( ethernet_mgmt.r_data         ),
            .s_axi_rresp    ( ethernet_mgmt.r_resp         ),
            .s_axi_rlast    ( ethernet_mgmt.r_last         ),
            .s_axi_rvalid   ( ethernet_mgmt.r_valid        ),
            .s_axi_rready   ( ethernet_mgmt.r_ready        ),

            .m_axi_awaddr   ( s_axi_ethernet_mgmt_awaddr   ),
            .m_axi_awlen    ( s_axi_ethernet_mgmt_awlen    ),
            .m_axi_awsize   ( s_axi_ethernet_mgmt_awsize   ),
            .m_axi_awburst  ( s_axi_ethernet_mgmt_awburst  ),
            .m_axi_awlock   ( s_axi_ethernet_mgmt_awlock   ),
            .m_axi_awcache  ( s_axi_ethernet_mgmt_awcache  ),
            .m_axi_awprot   ( s_axi_ethernet_mgmt_awprot   ),
            .m_axi_awregion ( s_axi_ethernet_mgmt_awregion ),
            .m_axi_awqos    ( s_axi_ethernet_mgmt_awqos    ),
            .m_axi_awvalid  ( s_axi_ethernet_mgmt_awvalid  ),
            .m_axi_awready  ( s_axi_ethernet_mgmt_awready  ),
            .m_axi_wdata    ( s_axi_ethernet_mgmt_wdata    ),
            .m_axi_wstrb    ( s_axi_ethernet_mgmt_wstrb    ),
            .m_axi_wlast    ( s_axi_ethernet_mgmt_wlast    ),
            .m_axi_wvalid   ( s_axi_ethernet_mgmt_wvalid   ),
            .m_axi_wready   ( s_axi_ethernet_mgmt_wready   ),
            .m_axi_bresp    ( s_axi_ethernet_mgmt_bresp    ),
            .m_axi_bvalid   ( s_axi_ethernet_mgmt_bvalid   ),
            .m_axi_bready   ( s_axi_ethernet_mgmt_bready   ),
            .m_axi_araddr   ( s_axi_ethernet_mgmt_araddr   ),
            .m_axi_arlen    ( s_axi_ethernet_mgmt_arlen    ),
            .m_axi_arsize   ( s_axi_ethernet_mgmt_arsize   ),
            .m_axi_arburst  ( s_axi_ethernet_mgmt_arburst  ),
            .m_axi_arlock   ( s_axi_ethernet_mgmt_arlock   ),
            .m_axi_arcache  ( s_axi_ethernet_mgmt_arcache  ),
            .m_axi_arprot   ( s_axi_ethernet_mgmt_arprot   ),
            .m_axi_arregion ( s_axi_ethernet_mgmt_arregion ),
            .m_axi_arqos    ( s_axi_ethernet_mgmt_arqos    ),
            .m_axi_arvalid  ( s_axi_ethernet_mgmt_arvalid  ),
            .m_axi_arready  ( s_axi_ethernet_mgmt_arready  ),
            .m_axi_rdata    ( s_axi_ethernet_mgmt_rdata    ),
            .m_axi_rresp    ( s_axi_ethernet_mgmt_rresp    ),
            .m_axi_rlast    ( s_axi_ethernet_mgmt_rlast    ),
            .m_axi_rvalid   ( s_axi_ethernet_mgmt_rvalid   ),
            .m_axi_rready   ( s_axi_ethernet_mgmt_rready   )
        );

        // Convert the full AXI ethernet MAC master into AXI lite
        logic [31:0] s_axi_lite_ethernet_mgmt_awaddr;
        logic        s_axi_lite_ethernet_mgmt_awvalid;
        logic        s_axi_lite_ethernet_mgmt_awready;
        logic [31:0] s_axi_lite_ethernet_mgmt_wdata;
        logic [3:0]  s_axi_lite_ethernet_mgmt_wstrb;
        logic        s_axi_lite_ethernet_mgmt_wvalid;
        logic        s_axi_lite_ethernet_mgmt_wready;
        logic [1:0]  s_axi_lite_ethernet_mgmt_bresp;
        logic        s_axi_lite_ethernet_mgmt_bvalid;
        logic        s_axi_lite_ethernet_mgmt_bready;
        logic [31:0] s_axi_lite_ethernet_mgmt_araddr;
        logic        s_axi_lite_ethernet_mgmt_arvalid;
        logic        s_axi_lite_ethernet_mgmt_arready;
        logic [31:0] s_axi_lite_ethernet_mgmt_rdata;
        logic [1:0]  s_axi_lite_ethernet_mgmt_rresp;
        logic        s_axi_lite_ethernet_mgmt_rvalid;
        logic        s_axi_lite_ethernet_mgmt_rready;

        xlnx_axi_lite_converter i_xlnx_axi_lite_converter_ethernet_mgmt (
            .aclk           ( clk_i                            ),
            .aresetn        ( rst_ni                           ),
            .s_axi_awaddr   ( s_axi_ethernet_mgmt_awaddr       ),
            .s_axi_awlen    ( s_axi_ethernet_mgmt_awlen        ),
            .s_axi_awsize   ( s_axi_ethernet_mgmt_awsize       ),
            .s_axi_awburst  ( s_axi_ethernet_mgmt_awburst      ),
            .s_axi_awlock   ( s_axi_ethernet_mgmt_awlock       ),
            .s_axi_awcache  ( s_axi_ethernet_mgmt_awcache      ),
            .s_axi_awprot   ( s_axi_ethernet_mgmt_awprot       ),
            .s_axi_awregion ( s_axi_ethernet_mgmt_awregion     ),
            .s_axi_awqos    ( s_axi_ethernet_mgmt_awqos        ),
            .s_axi_awvalid  ( s_axi_ethernet_mgmt_awvalid      ),
            .s_axi_awready  ( s_axi_ethernet_mgmt_awready      ),
            .s_axi_wdata    ( s_axi_ethernet_mgmt_wdata        ),
            .s_axi_wstrb    ( s_axi_ethernet_mgmt_wstrb        ),
            .s_axi_wlast    ( s_axi_ethernet_mgmt_wlast        ),
            .s_axi_wvalid   ( s_axi_ethernet_mgmt_wvalid       ),
            .s_axi_wready   ( s_axi_ethernet_mgmt_wready       ),
            .s_axi_bresp    ( s_axi_ethernet_mgmt_bresp        ),
            .s_axi_bvalid   ( s_axi_ethernet_mgmt_bvalid       ),
            .s_axi_bready   ( s_axi_ethernet_mgmt_bready       ),
            .s_axi_araddr   ( s_axi_ethernet_mgmt_araddr       ),
            .s_axi_arlen    ( s_axi_ethernet_mgmt_arlen        ),
            .s_axi_arsize   ( s_axi_ethernet_mgmt_arsize       ),
            .s_axi_arburst  ( s_axi_ethernet_mgmt_arburst      ),
            .s_axi_arlock   ( s_axi_ethernet_mgmt_arlock       ),
            .s_axi_arcache  ( s_axi_ethernet_mgmt_arcache      ),
            .s_axi_arprot   ( s_axi_ethernet_mgmt_arprot       ),
            .s_axi_arregion ( s_axi_ethernet_mgmt_arregion     ),
            .s_axi_arqos    ( s_axi_ethernet_mgmt_arqos        ),
            .s_axi_arvalid  ( s_axi_ethernet_mgmt_arvalid      ),
            .s_axi_arready  ( s_axi_ethernet_mgmt_arready      ),
            .s_axi_rdata    ( s_axi_ethernet_mgmt_rdata        ),
            .s_axi_rresp    ( s_axi_ethernet_mgmt_rresp        ),
            .s_axi_rlast    ( s_axi_ethernet_mgmt_rlast        ),
            .s_axi_rvalid   ( s_axi_ethernet_mgmt_rvalid       ),
            .s_axi_rready   ( s_axi_ethernet_mgmt_rready       ),

            .m_axi_awaddr   ( s_axi_lite_ethernet_mgmt_awaddr  ),
            .m_axi_awprot   ( /* NC */                         ),
            .m_axi_awvalid  ( s_axi_lite_ethernet_mgmt_awvalid ),
            .m_axi_awready  ( s_axi_lite_ethernet_mgmt_awready ),
            .m_axi_wdata    ( s_axi_lite_ethernet_mgmt_wdata   ),
            .m_axi_wstrb    ( s_axi_lite_ethernet_mgmt_wstrb   ),
            .m_axi_wvalid   ( s_axi_lite_ethernet_mgmt_wvalid  ),
            .m_axi_wready   ( s_axi_lite_ethernet_mgmt_wready  ),
            .m_axi_bresp    ( s_axi_lite_ethernet_mgmt_bresp   ),
            .m_axi_bvalid   ( s_axi_lite_ethernet_mgmt_bvalid  ),
            .m_axi_bready   ( s_axi_lite_ethernet_mgmt_bready  ),
            .m_axi_araddr   ( s_axi_lite_ethernet_mgmt_araddr  ),
            .m_axi_arprot   ( /* NC */                         ),
            .m_axi_arvalid  ( s_axi_lite_ethernet_mgmt_arvalid ),
            .m_axi_arready  ( s_axi_lite_ethernet_mgmt_arready ),
            .m_axi_rdata    ( s_axi_lite_ethernet_mgmt_rdata   ),
            .m_axi_rresp    ( s_axi_lite_ethernet_mgmt_rresp   ),
            .m_axi_rvalid   ( s_axi_lite_ethernet_mgmt_rvalid  ),
            .m_axi_rready   ( s_axi_lite_ethernet_mgmt_rready  )
        );

        // XXX The mdio signals from the MAC are not connected within the blackbox
        // axi_ethernet IP. The reason is unclear, but we are working on a fix.
        // Ethernet can work without it as the Phy will autonegotiate gigabit.

        xlnx_axi_ethernet i_xlnx_axi_ethernet_mac (
            .s_axi_lite_resetn      ( rst_ni                            ),
            .s_axi_lite_clk         ( clk_i                             ),
            // mac_irq isn't listed in the documentation. Perhaps it is
            // redundant with the "interrupt" wire?
            .mac_irq                ( /* NC */                          ),
            .axis_clk               ( clk_i                             ),
            .axi_txd_arstn          ( fifo_mm2s_prmry_reset_out_n       ),
            .axi_txc_arstn          ( fifo_mm2s_cntrl_reset_out_n       ),
            .axi_rxd_arstn          ( fifo_s2mm_prmry_reset_out_n       ),
            .axi_rxs_arstn          ( rst_ni                            ),
            .interrupt              ( irq_sources[2]                    ),
            .gtx_clk                ( phy_tx_clk_i                      ),
            .phy_rst_n              ( eth_rst_n                         ),
            .ref_clk                ( clk_200MHz_i                      ),
            // These clock outputs don't seem to be needed
            .gtx_clk90_out          ( /* NC */                          ),
            .gtx_clk_out            ( /* NC */                          ),
            .s_axi_araddr           ( s_axi_lite_ethernet_mgmt_araddr   ),
            .s_axi_arready          ( s_axi_lite_ethernet_mgmt_arready  ),
            .s_axi_arvalid          ( s_axi_lite_ethernet_mgmt_arvalid  ),
            .s_axi_awaddr           ( s_axi_lite_ethernet_mgmt_awaddr   ),
            .s_axi_awready          ( s_axi_lite_ethernet_mgmt_awready  ),
            .s_axi_awvalid          ( s_axi_lite_ethernet_mgmt_awvalid  ),
            .s_axi_bready           ( s_axi_lite_ethernet_mgmt_bready   ),
            .s_axi_bresp            ( s_axi_lite_ethernet_mgmt_bresp    ),
            .s_axi_bvalid           ( s_axi_lite_ethernet_mgmt_bvalid   ),
            .s_axi_rdata            ( s_axi_lite_ethernet_mgmt_rdata    ),
            .s_axi_rready           ( s_axi_lite_ethernet_mgmt_rready   ),
            .s_axi_rresp            ( s_axi_lite_ethernet_mgmt_rresp    ),
            .s_axi_rvalid           ( s_axi_lite_ethernet_mgmt_rvalid   ),
            .s_axi_wdata            ( s_axi_lite_ethernet_mgmt_wdata    ),
            .s_axi_wready           ( s_axi_lite_ethernet_mgmt_wready   ),
            .s_axi_wstrb            ( s_axi_lite_ethernet_mgmt_wstrb    ),
            .s_axi_wvalid           ( s_axi_lite_ethernet_mgmt_wvalid   ),
            .s_axis_txc_tdata       ( fifo_axi_str_txc_tdata            ),
            .s_axis_txc_tkeep       ( fifo_axi_str_txc_tkeep            ),
            .s_axis_txc_tlast       ( fifo_axi_str_txc_tlast            ),
            .s_axis_txc_tready      ( fifo_axi_str_txc_tready           ),
            .s_axis_txc_tvalid      ( fifo_axi_str_txc_tvalid           ),
            .s_axis_txd_tdata       ( fifo_axi_str_txd_tdata            ),
            .s_axis_txd_tkeep       ( fifo_axi_str_txd_tkeep            ),
            .s_axis_txd_tlast       ( fifo_axi_str_txd_tlast            ),
            .s_axis_txd_tready      ( fifo_axi_str_txd_tready           ),
            .s_axis_txd_tvalid      ( fifo_axi_str_txd_tvalid           ),
            .m_axis_rxd_tdata       ( fifo_axi_str_rxd_tdata            ),
            .m_axis_rxd_tkeep       ( fifo_axi_str_rxd_tkeep            ),
            .m_axis_rxd_tlast       ( fifo_axi_str_rxd_tlast            ),
            .m_axis_rxd_tready      ( fifo_axi_str_rxd_tready           ),
            .m_axis_rxd_tvalid      ( fifo_axi_str_rxd_tvalid           ),
            // The specification gives the case of connecting to the FIFO
            // as an example, specifying these connections
            .m_axis_rxs_tdata       ( /* NC */                          ),
            .m_axis_rxs_tkeep       ( /* NC */                          ),
            .m_axis_rxs_tlast       ( /* NC */                          ),
            .m_axis_rxs_tready      ( 1'b1                              ),
            .m_axis_rxs_tvalid      ( /* NC */                          ),
            .rgmii_rd               ( eth_rxd                           ),
            .rgmii_rx_ctl           ( eth_rxctl                         ),
            .rgmii_rxc              ( eth_rxck                          ),
            .rgmii_td               ( eth_txd                           ),
            .rgmii_tx_ctl           ( eth_txctl                         ),
            .rgmii_txc              ( eth_txck                          ),
            .mdio_mdc               ( eth_mdc                           ),
            .mdio_mdio_i            ( eth_mdio_i                        ),
            .mdio_mdio_o            ( eth_mdio_o                        ),
            .mdio_mdio_t            ( eth_mdio_oe                       )
        );
    end else begin
        // Tie off signals with no separate ethernet management interface
        assign irq_sources [7] = 1'b0;
        assign ethernet_mgmt.aw_ready = 1'b1;
        assign ethernet_mgmt.ar_ready = 1'b1;
        assign ethernet_mgmt.w_ready = 1'b1;

        assign ethernet_mgmt.b_valid = ethernet_mgmt.aw_valid;
        assign ethernet_mgmt.b_id = ethernet_mgmt.aw_id;
        assign ethernet_mgmt.b_resp = axi_pkg::RESP_SLVERR;
        assign ethernet_mgmt.b_user = '0;

        assign ethernet_mgmt.r_valid = ethernet_mgmt.ar_valid;
        assign ethernet_mgmt.r_resp = axi_pkg::RESP_SLVERR;
        assign ethernet_mgmt.r_data = 'hdeadbeef;
        assign ethernet_mgmt.r_last = 1'b1;
    end

    if (InclLowriscEthernet) begin : gen_lowrisc_ethernet
        logic                    clk_200_int, clk_rgmii, clk_rgmii_quad;
        logic                    eth_en, eth_we, eth_int_n, eth_pme_n;
        logic [AxiAddrWidth-1:0] eth_addr;
        logic [AxiDataWidth-1:0] eth_wrdata, eth_rdata;
        logic [AxiDataWidth/8-1:0] eth_be;

        axi2mem #(
            .AXI_ID_WIDTH   ( AxiIdWidth   ),
            .AXI_ADDR_WIDTH ( AxiAddrWidth ),
            .AXI_DATA_WIDTH ( AxiDataWidth ),
            .AXI_USER_WIDTH ( AxiUserWidth )
        ) i_axi2rom (
            .clk_i  ( clk_i         ),
            .rst_ni ( rst_ni        ),
            .slave  ( ethernet_data ),
            .req_o  ( eth_en        ),
            .we_o   ( eth_we        ),
            .addr_o ( eth_addr      ),
            .be_o   ( eth_be        ),
            .data_o ( eth_wrdata    ),
            .data_i ( eth_rdata     )
        );

        framing_top eth_rgmii (
           .msoc_clk(clk_i),
           .core_lsu_addr(eth_addr[14:0]),
           .core_lsu_wdata(eth_wrdata),
           .core_lsu_be(eth_be),
           .ce_d(eth_en),
           .we_d(eth_en & eth_we),
           .framing_sel(eth_en),
           .framing_rdata(eth_rdata),
           .rst_int(!rst_ni),
           .clk_int(phy_tx_clk_i), // 125 MHz in-phase
           .clk90_int(eth_clk_i),    // 125 MHz quadrature
           .clk_200_int(clk_200MHz_i),
           /*
            * Ethernet: 1000BASE-T RGMII
            */
           .phy_rx_clk(eth_rxck),
           .phy_rxd(eth_rxd),
           .phy_rx_ctl(eth_rxctl),
           .phy_tx_clk(eth_txck),
           .phy_txd(eth_txd),
           .phy_tx_ctl(eth_txctl),
           .phy_reset_n(eth_rst_n),
           .phy_int_n(eth_int_n),
           .phy_pme_n(eth_pme_n),
           .phy_mdc(eth_mdc),
           .phy_mdio_i(eth_mdio_i),
           .phy_mdio_o(eth_mdio_o),
           .phy_mdio_oe(~eth_mdio_oe),
           .eth_irq(irq_sources[2])
        );
    end

    // 5. GPIO
    assign gpio.b_user = 1'b0;
    assign gpio.r_user = 1'b0;

    if (InclGPIO) begin : gen_gpio

        logic [31:0] s_axi_gpio_awaddr;
        logic [7:0]  s_axi_gpio_awlen;
        logic [2:0]  s_axi_gpio_awsize;
        logic [1:0]  s_axi_gpio_awburst;
        logic [3:0]  s_axi_gpio_awcache;
        logic        s_axi_gpio_awvalid;
        logic        s_axi_gpio_awready;
        logic [31:0] s_axi_gpio_wdata;
        logic [3:0]  s_axi_gpio_wstrb;
        logic        s_axi_gpio_wvalid;
        logic        s_axi_gpio_wready;
        logic [1:0]  s_axi_gpio_bresp;
        logic        s_axi_gpio_bvalid;
        logic        s_axi_gpio_bready;
        logic [31:0] s_axi_gpio_araddr;
        logic [7:0]  s_axi_gpio_arlen;
        logic [2:0]  s_axi_gpio_arsize;
        logic [1:0]  s_axi_gpio_arburst;
        logic [3:0]  s_axi_gpio_arcache;
        logic        s_axi_gpio_arvalid;
        logic        s_axi_gpio_arready;
        logic [31:0] s_axi_gpio_rdata;
        logic [1:0]  s_axi_gpio_rresp;
        logic        s_axi_gpio_rlast;
        logic        s_axi_gpio_rvalid;
        logic        s_axi_gpio_rready;

        // system-bus is 64-bit, convert down to 32 bit
        xlnx_axi_dwidth_converter i_xlnx_axi_dwidth_converter_gpio (
            .s_axi_aclk     ( clk_i              ),
            .s_axi_aresetn  ( rst_ni             ),
            .s_axi_awid     ( gpio.aw_id         ),
            .s_axi_awaddr   ( gpio.aw_addr[31:0] ),
            .s_axi_awlen    ( gpio.aw_len        ),
            .s_axi_awsize   ( gpio.aw_size       ),
            .s_axi_awburst  ( gpio.aw_burst      ),
            .s_axi_awlock   ( gpio.aw_lock       ),
            .s_axi_awcache  ( gpio.aw_cache      ),
            .s_axi_awprot   ( gpio.aw_prot       ),
            .s_axi_awregion ( gpio.aw_region     ),
            .s_axi_awqos    ( gpio.aw_qos        ),
            .s_axi_awvalid  ( gpio.aw_valid      ),
            .s_axi_awready  ( gpio.aw_ready      ),
            .s_axi_wdata    ( gpio.w_data        ),
            .s_axi_wstrb    ( gpio.w_strb        ),
            .s_axi_wlast    ( gpio.w_last        ),
            .s_axi_wvalid   ( gpio.w_valid       ),
            .s_axi_wready   ( gpio.w_ready       ),
            .s_axi_bid      ( gpio.b_id          ),
            .s_axi_bresp    ( gpio.b_resp        ),
            .s_axi_bvalid   ( gpio.b_valid       ),
            .s_axi_bready   ( gpio.b_ready       ),
            .s_axi_arid     ( gpio.ar_id         ),
            .s_axi_araddr   ( gpio.ar_addr[31:0] ),
            .s_axi_arlen    ( gpio.ar_len        ),
            .s_axi_arsize   ( gpio.ar_size       ),
            .s_axi_arburst  ( gpio.ar_burst      ),
            .s_axi_arlock   ( gpio.ar_lock       ),
            .s_axi_arcache  ( gpio.ar_cache      ),
            .s_axi_arprot   ( gpio.ar_prot       ),
            .s_axi_arregion ( gpio.ar_region     ),
            .s_axi_arqos    ( gpio.ar_qos        ),
            .s_axi_arvalid  ( gpio.ar_valid      ),
            .s_axi_arready  ( gpio.ar_ready      ),
            .s_axi_rid      ( gpio.r_id          ),
            .s_axi_rdata    ( gpio.r_data        ),
            .s_axi_rresp    ( gpio.r_resp        ),
            .s_axi_rlast    ( gpio.r_last        ),
            .s_axi_rvalid   ( gpio.r_valid       ),
            .s_axi_rready   ( gpio.r_ready       ),

            .m_axi_awaddr   ( s_axi_gpio_awaddr  ),
            .m_axi_awlen    ( s_axi_gpio_awlen   ),
            .m_axi_awsize   ( s_axi_gpio_awsize  ),
            .m_axi_awburst  ( s_axi_gpio_awburst ),
            .m_axi_awlock   (                    ),
            .m_axi_awcache  ( s_axi_gpio_awcache ),
            .m_axi_awprot   (                    ),
            .m_axi_awregion (                    ),
            .m_axi_awqos    (                    ),
            .m_axi_awvalid  ( s_axi_gpio_awvalid ),
            .m_axi_awready  ( s_axi_gpio_awready ),
            .m_axi_wdata    ( s_axi_gpio_wdata   ),
            .m_axi_wstrb    ( s_axi_gpio_wstrb   ),
            .m_axi_wlast    (                    ),
            .m_axi_wvalid   ( s_axi_gpio_wvalid  ),
            .m_axi_wready   ( s_axi_gpio_wready  ),
            .m_axi_bresp    ( s_axi_gpio_bresp   ),
            .m_axi_bvalid   ( s_axi_gpio_bvalid  ),
            .m_axi_bready   ( s_axi_gpio_bready  ),
            .m_axi_araddr   ( s_axi_gpio_araddr  ),
            .m_axi_arlen    ( s_axi_gpio_arlen   ),
            .m_axi_arsize   ( s_axi_gpio_arsize  ),
            .m_axi_arburst  ( s_axi_gpio_arburst ),
            .m_axi_arlock   (                    ),
            .m_axi_arcache  ( s_axi_gpio_arcache ),
            .m_axi_arprot   (                    ),
            .m_axi_arregion (                    ),
            .m_axi_arqos    (                    ),
            .m_axi_arvalid  ( s_axi_gpio_arvalid ),
            .m_axi_arready  ( s_axi_gpio_arready ),
            .m_axi_rdata    ( s_axi_gpio_rdata   ),
            .m_axi_rresp    ( s_axi_gpio_rresp   ),
            .m_axi_rlast    ( s_axi_gpio_rlast   ),
            .m_axi_rvalid   ( s_axi_gpio_rvalid  ),
            .m_axi_rready   ( s_axi_gpio_rready  )
        );

        xlnx_axi_gpio i_xlnx_axi_gpio (
            .s_axi_aclk    ( clk_i                  ),
            .s_axi_aresetn ( rst_ni                 ),
            .s_axi_awaddr  ( s_axi_gpio_awaddr[8:0] ),
            .s_axi_awvalid ( s_axi_gpio_awvalid     ),
            .s_axi_awready ( s_axi_gpio_awready     ),
            .s_axi_wdata   ( s_axi_gpio_wdata       ),
            .s_axi_wstrb   ( s_axi_gpio_wstrb       ),
            .s_axi_wvalid  ( s_axi_gpio_wvalid      ),
            .s_axi_wready  ( s_axi_gpio_wready      ),
            .s_axi_bresp   ( s_axi_gpio_bresp       ),
            .s_axi_bvalid  ( s_axi_gpio_bvalid      ),
            .s_axi_bready  ( s_axi_gpio_bready      ),
            .s_axi_araddr  ( s_axi_gpio_araddr[8:0] ),
            .s_axi_arvalid ( s_axi_gpio_arvalid     ),
            .s_axi_arready ( s_axi_gpio_arready     ),
            .s_axi_rdata   ( s_axi_gpio_rdata       ),
            .s_axi_rresp   ( s_axi_gpio_rresp       ),
            .s_axi_rvalid  ( s_axi_gpio_rvalid      ),
            .s_axi_rready  ( s_axi_gpio_rready      ),
            .gpio_io_i     ( '0                     ),
            .gpio_io_o     ( leds_o                 ),
            .gpio_io_t     (                        ),
            .gpio2_io_i    ( dip_switches_i         )
        );

        assign s_axi_gpio_rlast = 1'b1;

    end

    // 6. Timer
    if (InclTimer) begin : gen_timer
        logic         timer_penable;
        logic         timer_pwrite;
        logic [31:0]  timer_paddr;
        logic         timer_psel;
        logic [31:0]  timer_pwdata;
        logic [31:0]  timer_prdata;
        logic         timer_pready;
        logic         timer_pslverr;

        axi2apb_64_32 #(
            .AXI4_ADDRESS_WIDTH ( AxiAddrWidth ),
            .AXI4_RDATA_WIDTH   ( AxiDataWidth ),
            .AXI4_WDATA_WIDTH   ( AxiDataWidth ),
            .AXI4_ID_WIDTH      ( AxiIdWidth   ),
            .AXI4_USER_WIDTH    ( AxiUserWidth ),
            .BUFF_DEPTH_SLAVE   ( 2            ),
            .APB_ADDR_WIDTH     ( 32           )
        ) i_axi2apb_64_32_timer (
            .ACLK      ( clk_i           ),
            .ARESETn   ( rst_ni          ),
            .test_en_i ( 1'b0            ),
            .AWID_i    ( timer.aw_id     ),
            .AWADDR_i  ( timer.aw_addr   ),
            .AWLEN_i   ( timer.aw_len    ),
            .AWSIZE_i  ( timer.aw_size   ),
            .AWBURST_i ( timer.aw_burst  ),
            .AWLOCK_i  ( timer.aw_lock   ),
            .AWCACHE_i ( timer.aw_cache  ),
            .AWPROT_i  ( timer.aw_prot   ),
            .AWREGION_i( timer.aw_region ),
            .AWUSER_i  ( timer.aw_user   ),
            .AWQOS_i   ( timer.aw_qos    ),
            .AWVALID_i ( timer.aw_valid  ),
            .AWREADY_o ( timer.aw_ready  ),
            .WDATA_i   ( timer.w_data    ),
            .WSTRB_i   ( timer.w_strb    ),
            .WLAST_i   ( timer.w_last    ),
            .WUSER_i   ( timer.w_user    ),
            .WVALID_i  ( timer.w_valid   ),
            .WREADY_o  ( timer.w_ready   ),
            .BID_o     ( timer.b_id      ),
            .BRESP_o   ( timer.b_resp    ),
            .BVALID_o  ( timer.b_valid   ),
            .BUSER_o   ( timer.b_user    ),
            .BREADY_i  ( timer.b_ready   ),
            .ARID_i    ( timer.ar_id     ),
            .ARADDR_i  ( timer.ar_addr   ),
            .ARLEN_i   ( timer.ar_len    ),
            .ARSIZE_i  ( timer.ar_size   ),
            .ARBURST_i ( timer.ar_burst  ),
            .ARLOCK_i  ( timer.ar_lock   ),
            .ARCACHE_i ( timer.ar_cache  ),
            .ARPROT_i  ( timer.ar_prot   ),
            .ARREGION_i( timer.ar_region ),
            .ARUSER_i  ( timer.ar_user   ),
            .ARQOS_i   ( timer.ar_qos    ),
            .ARVALID_i ( timer.ar_valid  ),
            .ARREADY_o ( timer.ar_ready  ),
            .RID_o     ( timer.r_id      ),
            .RDATA_o   ( timer.r_data    ),
            .RRESP_o   ( timer.r_resp    ),
            .RLAST_o   ( timer.r_last    ),
            .RUSER_o   ( timer.r_user    ),
            .RVALID_o  ( timer.r_valid   ),
            .RREADY_i  ( timer.r_ready   ),
            .PENABLE   ( timer_penable   ),
            .PWRITE    ( timer_pwrite    ),
            .PADDR     ( timer_paddr     ),
            .PSEL      ( timer_psel      ),
            .PWDATA    ( timer_pwdata    ),
            .PRDATA    ( timer_prdata    ),
            .PREADY    ( timer_pready    ),
            .PSLVERR   ( timer_pslverr   )
        );

        apb_timer #(
                .APB_ADDR_WIDTH ( 32 ),
                .TIMER_CNT      ( 2  )
        ) i_timer (
            .HCLK    ( clk_i            ),
            .HRESETn ( rst_ni           ),
            .PSEL    ( timer_psel       ),
            .PENABLE ( timer_penable    ),
            .PWRITE  ( timer_pwrite     ),
            .PADDR   ( timer_paddr      ),
            .PWDATA  ( timer_pwdata     ),
            .PRDATA  ( timer_prdata     ),
            .PREADY  ( timer_pready     ),
            .PSLVERR ( timer_pslverr    ),
            .irq_o   ( irq_sources[6:3] )
        );
    end
endmodule
